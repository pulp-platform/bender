module leaf;
endmodule
