module unused_top;
    unused_leaf u_unused_leaf();
endmodule
