module core;
    leaf u_leaf();
endmodule
