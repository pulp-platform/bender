module unused_leaf;
endmodule
