module broken(;
endmodule
