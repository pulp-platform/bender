// Module with a named end label to test that `endmodule : name` is also renamed.
module named_end;
endmodule : named_end
